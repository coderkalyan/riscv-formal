../../../discrete_rvfi_monitor.vh